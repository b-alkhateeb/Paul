module dff(x,y,z);

endmodule